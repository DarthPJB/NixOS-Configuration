* Simple Voltage Divider Circuit
V1 in 0 5
R1 in out 1k
R2 out 0 1k
.dc
.print dc V(out)
.end
