* Simple Voltage Divider Circuit
V1 1 0 DC 5V
R1 1 out 1k
R2 out 0 1k
.PRINT DC V(out)
.DC
.end
